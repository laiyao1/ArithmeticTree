module main(a,b,s,cout);
input [63:0] a,b;
output [63:0] s;
output cout;
wire p39_36,g43_43,p17_17,g15_8,p26_23,g28_23,p27_26,p9_9,g56_55,g5_0,p40_33,g31_22,g4_4,g63_63,p3_3,g35_33,c41,p0_0,p45_45,p14_8,g6_6,g41_33,c6,c53,g40_36,g25_25,c63,c54,p13_13,g26_23,p22_22,g32_23,p26_26,g51_50,p58_41,p8_8,g19_19,g55_55,c2,p39_33,g57_55,g6_0,g15_15,c29,g39_36,p29_29,g3_0,p55_55,c17,p57_55,g0_0,g3_3,g34_33,p56_55,g22_22,c36,g49_42,g44_42,p46_42,c40,p35_33,p48_48,p15_8,c51,p41_23,p29_23,g34_34,p49_49,g9_7,p33_33,g16_0,p56_42,c30,g60_42,c60,g37_33,g58_41,g57_42,p51_42,c3,p55_23,c15,p25_23,p24_24,c24,g1_1,g9_9,c19,p56_56,c28,p18_18,g41_23,p5_5,c58,c55,g58_42,g10_8,c46,g16_16,g35_35,g52_52,c11,g62_62,p32_23,p2_2,g37_36,p39_39,g49_0,p6_6,g45_45,p44_42,p42_42,p27_23,g31_31,g59_59,g10_10,g7_0,p60_60,g26_26,p37_33,p35_35,p36_36,g47_42,p10_10,p58_58,p57_42,c31,g28_28,g11_11,g12_12,p47_42,g1_0,g30_23,g42_42,c39,p4_4,p53_53,c57,c34,c61,p28_23,c38,p30_30,g13_13,p48_42,g29_23,c10,p38_36,g37_37,p1_1,g58_58,g48_42,p49_42,p41_41,p16_16,g18_18,p54_23,c14,g14_14,g45_42,g36_36,c48,g15_0,p58_42,c16,p12_8,g33_33,g2_0,g8_8,p51_51,p15_15,g13_8,p47_47,p27_27,p40_40,g18_0,g21_21,g46_42,g32_32,g7_7,c12,c21,g12_8,g20_20,g41_41,g9_8,g21_0,p50_50,p38_33,c22,p9_8,p41_33,g40_33,p59_59,g23_23,c37,g61_61,c49,c27,c13,g40_0,g43_42,g60_60,p60_42,p63_63,g49_49,p20_20,c50,p10_8,c1,p61_61,g39_39,p28_28,p37_36,p14_14,c59,g46_46,g56_42,g54_23,g59_42,c7,p34_34,g51_51,p51_50,p46_46,c47,c43,p30_23,p52_52,p11_8,g14_8,c4,p43_42,p59_42,c5,g62_0,c18,g27_23,c25,p31_31,g27_26,p61_42,g40_40,p54_54,g2_2,g54_42,p57_57,p12_12,p31_22,c8,p34_33,g17_0,p32_32,c9,p25_25,c33,p11_11,g11_8,g4_0,c20,p44_44,g52_42,g24_24,p21_21,g61_42,g44_44,g17_17,g24_23,g38_38,c44,c52,g27_27,g5_5,g53_53,p38_38,p31_23,g30_30,g39_33,g54_54,p23_23,g53_42,p19_19,g35_0,c32,g31_23,g50_50,c23,p53_42,p7_7,p9_7,g29_29,g48_48,p40_36,g19_0,p52_42,c45,p62_62,p45_42,g41_0,c0,p13_8,g57_57,c26,c35,c56,c42,g55_23,g20_0,c62,g38_33,g56_56,g32_0,g47_47,p37_37,g38_36,g25_23,p24_23,g22_0,p54_42,p43_43,g61_0,g51_42;

assign p0_0 = a[0] ^ b[0];
assign g0_0 = a[0] & b[0];
assign p1_1 = a[1] ^ b[1];
assign g1_1 = a[1] & b[1];
assign p2_2 = a[2] ^ b[2];
assign g2_2 = a[2] & b[2];
assign p3_3 = a[3] ^ b[3];
assign g3_3 = a[3] & b[3];
assign p4_4 = a[4] ^ b[4];
assign g4_4 = a[4] & b[4];
assign p5_5 = a[5] ^ b[5];
assign g5_5 = a[5] & b[5];
assign p6_6 = a[6] ^ b[6];
assign g6_6 = a[6] & b[6];
assign p7_7 = a[7] ^ b[7];
assign g7_7 = a[7] & b[7];
assign p8_8 = a[8] ^ b[8];
assign g8_8 = a[8] & b[8];
assign p9_9 = a[9] ^ b[9];
assign g9_9 = a[9] & b[9];
assign p10_10 = a[10] ^ b[10];
assign g10_10 = a[10] & b[10];
assign p11_11 = a[11] ^ b[11];
assign g11_11 = a[11] & b[11];
assign p12_12 = a[12] ^ b[12];
assign g12_12 = a[12] & b[12];
assign p13_13 = a[13] ^ b[13];
assign g13_13 = a[13] & b[13];
assign p14_14 = a[14] ^ b[14];
assign g14_14 = a[14] & b[14];
assign p15_15 = a[15] ^ b[15];
assign g15_15 = a[15] & b[15];
assign p16_16 = a[16] ^ b[16];
assign g16_16 = a[16] & b[16];
assign p17_17 = a[17] ^ b[17];
assign g17_17 = a[17] & b[17];
assign p18_18 = a[18] ^ b[18];
assign g18_18 = a[18] & b[18];
assign p19_19 = a[19] ^ b[19];
assign g19_19 = a[19] & b[19];
assign p20_20 = a[20] ^ b[20];
assign g20_20 = a[20] & b[20];
assign p21_21 = a[21] ^ b[21];
assign g21_21 = a[21] & b[21];
assign p22_22 = a[22] ^ b[22];
assign g22_22 = a[22] & b[22];
assign p23_23 = a[23] ^ b[23];
assign g23_23 = a[23] & b[23];
assign p24_24 = a[24] ^ b[24];
assign g24_24 = a[24] & b[24];
assign p25_25 = a[25] ^ b[25];
assign g25_25 = a[25] & b[25];
assign p26_26 = a[26] ^ b[26];
assign g26_26 = a[26] & b[26];
assign p27_27 = a[27] ^ b[27];
assign g27_27 = a[27] & b[27];
assign p28_28 = a[28] ^ b[28];
assign g28_28 = a[28] & b[28];
assign p29_29 = a[29] ^ b[29];
assign g29_29 = a[29] & b[29];
assign p30_30 = a[30] ^ b[30];
assign g30_30 = a[30] & b[30];
assign p31_31 = a[31] ^ b[31];
assign g31_31 = a[31] & b[31];
assign p32_32 = a[32] ^ b[32];
assign g32_32 = a[32] & b[32];
assign p33_33 = a[33] ^ b[33];
assign g33_33 = a[33] & b[33];
assign p34_34 = a[34] ^ b[34];
assign g34_34 = a[34] & b[34];
assign p35_35 = a[35] ^ b[35];
assign g35_35 = a[35] & b[35];
assign p36_36 = a[36] ^ b[36];
assign g36_36 = a[36] & b[36];
assign p37_37 = a[37] ^ b[37];
assign g37_37 = a[37] & b[37];
assign p38_38 = a[38] ^ b[38];
assign g38_38 = a[38] & b[38];
assign p39_39 = a[39] ^ b[39];
assign g39_39 = a[39] & b[39];
assign p40_40 = a[40] ^ b[40];
assign g40_40 = a[40] & b[40];
assign p41_41 = a[41] ^ b[41];
assign g41_41 = a[41] & b[41];
assign p42_42 = a[42] ^ b[42];
assign g42_42 = a[42] & b[42];
assign p43_43 = a[43] ^ b[43];
assign g43_43 = a[43] & b[43];
assign p44_44 = a[44] ^ b[44];
assign g44_44 = a[44] & b[44];
assign p45_45 = a[45] ^ b[45];
assign g45_45 = a[45] & b[45];
assign p46_46 = a[46] ^ b[46];
assign g46_46 = a[46] & b[46];
assign p47_47 = a[47] ^ b[47];
assign g47_47 = a[47] & b[47];
assign p48_48 = a[48] ^ b[48];
assign g48_48 = a[48] & b[48];
assign p49_49 = a[49] ^ b[49];
assign g49_49 = a[49] & b[49];
assign p50_50 = a[50] ^ b[50];
assign g50_50 = a[50] & b[50];
assign p51_51 = a[51] ^ b[51];
assign g51_51 = a[51] & b[51];
assign p52_52 = a[52] ^ b[52];
assign g52_52 = a[52] & b[52];
assign p53_53 = a[53] ^ b[53];
assign g53_53 = a[53] & b[53];
assign p54_54 = a[54] ^ b[54];
assign g54_54 = a[54] & b[54];
assign p55_55 = a[55] ^ b[55];
assign g55_55 = a[55] & b[55];
assign p56_56 = a[56] ^ b[56];
assign g56_56 = a[56] & b[56];
assign p57_57 = a[57] ^ b[57];
assign g57_57 = a[57] & b[57];
assign p58_58 = a[58] ^ b[58];
assign g58_58 = a[58] & b[58];
assign p59_59 = a[59] ^ b[59];
assign g59_59 = a[59] & b[59];
assign p60_60 = a[60] ^ b[60];
assign g60_60 = a[60] & b[60];
assign p61_61 = a[61] ^ b[61];
assign g61_61 = a[61] & b[61];
assign p62_62 = a[62] ^ b[62];
assign g62_62 = a[62] & b[62];
assign p63_63 = a[63] ^ b[63];
assign g63_63 = a[63] & b[63];
assign g1_0 = c1;
assign g2_0 = c2;
assign g3_0 = c3;
assign g4_0 = c4;
assign g5_0 = c5;
assign g6_0 = c6;
assign g7_0 = c7;
assign g8_0 = c8;
assign g9_0 = c9;
assign g10_0 = c10;
assign g11_0 = c11;
assign g12_0 = c12;
assign g13_0 = c13;
assign g14_0 = c14;
assign g15_0 = c15;
assign g16_0 = c16;
assign g17_0 = c17;
assign g18_0 = c18;
assign g19_0 = c19;
assign g20_0 = c20;
assign g21_0 = c21;
assign g22_0 = c22;
assign g23_0 = c23;
assign g24_0 = c24;
assign g25_0 = c25;
assign g26_0 = c26;
assign g27_0 = c27;
assign g28_0 = c28;
assign g29_0 = c29;
assign g30_0 = c30;
assign g31_0 = c31;
assign g32_0 = c32;
assign g33_0 = c33;
assign g34_0 = c34;
assign g35_0 = c35;
assign g36_0 = c36;
assign g37_0 = c37;
assign g38_0 = c38;
assign g39_0 = c39;
assign g40_0 = c40;
assign g41_0 = c41;
assign g42_0 = c42;
assign g43_0 = c43;
assign g44_0 = c44;
assign g45_0 = c45;
assign g46_0 = c46;
assign g47_0 = c47;
assign g48_0 = c48;
assign g49_0 = c49;
assign g50_0 = c50;
assign g51_0 = c51;
assign g52_0 = c52;
assign g53_0 = c53;
assign g54_0 = c54;
assign g55_0 = c55;
assign g56_0 = c56;
assign g57_0 = c57;
assign g58_0 = c58;
assign g59_0 = c59;
assign g60_0 = c60;
assign g61_0 = c61;
assign g62_0 = c62;
assign g63_0 = c63;
GREY grey63(g63_63, p63_63, g62_0, c63);
GREY grey62(g62_62, p62_62, g61_0, c62);
BLACK black61_42(g61_61, p61_61, g60_42, p60_42, g61_42, p61_42);
GREY grey61(g61_42, p61_42, g41_0, c61);
BLACK black60_42(g60_60, p60_60, g59_42, p59_42, g60_42, p60_42);
GREY grey60(g60_42, p60_42, g41_0, c60);
BLACK black59_42(g59_59, p59_59, g58_42, p58_42, g59_42, p59_42);
GREY grey59(g59_42, p59_42, g41_0, c59);
BLACK black58_42(g58_58, p58_58, g57_42, p57_42, g58_42, p58_42);
BLACK black58_41(g58_42, p58_42, g41_41, p41_41, g58_41, p58_41);
GREY grey58(g58_41, p58_41, g40_0, c58);
BLACK black57_55(g57_57, p57_57, g56_55, p56_55, g57_55, p57_55);
BLACK black57_42(g57_55, p57_55, g54_42, p54_42, g57_42, p57_42);
GREY grey57(g57_42, p57_42, g41_0, c57);
BLACK black56_55(g56_56, p56_56, g55_55, p55_55, g56_55, p56_55);
BLACK black56_42(g56_55, p56_55, g54_42, p54_42, g56_42, p56_42);
GREY grey56(g56_42, p56_42, g41_0, c56);
BLACK black55_23(g55_55, p55_55, g54_23, p54_23, g55_23, p55_23);
GREY grey55(g55_23, p55_23, g22_0, c55);
BLACK black54_42(g54_54, p54_54, g53_42, p53_42, g54_42, p54_42);
BLACK black54_23(g54_42, p54_42, g41_23, p41_23, g54_23, p54_23);
GREY grey54(g54_23, p54_23, g22_0, c54);
BLACK black53_42(g53_53, p53_53, g52_42, p52_42, g53_42, p53_42);
GREY grey53(g53_42, p53_42, g41_0, c53);
BLACK black52_42(g52_52, p52_52, g51_42, p51_42, g52_42, p52_42);
GREY grey52(g52_42, p52_42, g41_0, c52);
BLACK black51_50(g51_51, p51_51, g50_50, p50_50, g51_50, p51_50);
BLACK black51_42(g51_50, p51_50, g49_42, p49_42, g51_42, p51_42);
GREY grey51(g51_42, p51_42, g41_0, c51);
GREY grey50(g50_50, p50_50, g49_0, c50);
BLACK black49_42(g49_49, p49_49, g48_42, p48_42, g49_42, p49_42);
GREY grey49(g49_42, p49_42, g41_0, c49);
BLACK black48_42(g48_48, p48_48, g47_42, p47_42, g48_42, p48_42);
GREY grey48(g48_42, p48_42, g41_0, c48);
BLACK black47_42(g47_47, p47_47, g46_42, p46_42, g47_42, p47_42);
GREY grey47(g47_42, p47_42, g41_0, c47);
BLACK black46_42(g46_46, p46_46, g45_42, p45_42, g46_42, p46_42);
GREY grey46(g46_42, p46_42, g41_0, c46);
BLACK black45_42(g45_45, p45_45, g44_42, p44_42, g45_42, p45_42);
GREY grey45(g45_42, p45_42, g41_0, c45);
BLACK black44_42(g44_44, p44_44, g43_42, p43_42, g44_42, p44_42);
GREY grey44(g44_42, p44_42, g41_0, c44);
BLACK black43_42(g43_43, p43_43, g42_42, p42_42, g43_42, p43_42);
GREY grey43(g43_42, p43_42, g41_0, c43);
GREY grey42(g42_42, p42_42, g41_0, c42);
BLACK black41_33(g41_41, p41_41, g40_33, p40_33, g41_33, p41_33);
BLACK black41_23(g41_33, p41_33, g32_23, p32_23, g41_23, p41_23);
GREY grey41(g41_23, p41_23, g22_0, c41);
BLACK black40_36(g40_40, p40_40, g39_36, p39_36, g40_36, p40_36);
BLACK black40_33(g40_36, p40_36, g35_33, p35_33, g40_33, p40_33);
GREY grey40(g40_33, p40_33, g32_0, c40);
BLACK black39_36(g39_39, p39_39, g38_36, p38_36, g39_36, p39_36);
BLACK black39_33(g39_36, p39_36, g35_33, p35_33, g39_33, p39_33);
GREY grey39(g39_33, p39_33, g32_0, c39);
BLACK black38_36(g38_38, p38_38, g37_36, p37_36, g38_36, p38_36);
BLACK black38_33(g38_36, p38_36, g35_33, p35_33, g38_33, p38_33);
GREY grey38(g38_33, p38_33, g32_0, c38);
BLACK black37_36(g37_37, p37_37, g36_36, p36_36, g37_36, p37_36);
BLACK black37_33(g37_36, p37_36, g35_33, p35_33, g37_33, p37_33);
GREY grey37(g37_33, p37_33, g32_0, c37);
GREY grey36(g36_36, p36_36, g35_0, c36);
BLACK black35_33(g35_35, p35_35, g34_33, p34_33, g35_33, p35_33);
GREY grey35(g35_33, p35_33, g32_0, c35);
BLACK black34_33(g34_34, p34_34, g33_33, p33_33, g34_33, p34_33);
GREY grey34(g34_33, p34_33, g32_0, c34);
GREY grey33(g33_33, p33_33, g32_0, c33);
BLACK black32_23(g32_32, p32_32, g31_23, p31_23, g32_23, p32_23);
GREY grey32(g32_23, p32_23, g22_0, c32);
BLACK black31_23(g31_31, p31_31, g30_23, p30_23, g31_23, p31_23);
BLACK black31_22(g31_23, p31_23, g22_22, p22_22, g31_22, p31_22);
GREY grey31(g31_22, p31_22, g21_0, c31);
BLACK black30_23(g30_30, p30_30, g29_23, p29_23, g30_23, p30_23);
GREY grey30(g30_23, p30_23, g22_0, c30);
BLACK black29_23(g29_29, p29_29, g28_23, p28_23, g29_23, p29_23);
GREY grey29(g29_23, p29_23, g22_0, c29);
BLACK black28_23(g28_28, p28_28, g27_23, p27_23, g28_23, p28_23);
GREY grey28(g28_23, p28_23, g22_0, c28);
BLACK black27_26(g27_27, p27_27, g26_26, p26_26, g27_26, p27_26);
BLACK black27_23(g27_26, p27_26, g25_23, p25_23, g27_23, p27_23);
GREY grey27(g27_23, p27_23, g22_0, c27);
BLACK black26_23(g26_26, p26_26, g25_23, p25_23, g26_23, p26_23);
GREY grey26(g26_23, p26_23, g22_0, c26);
BLACK black25_23(g25_25, p25_25, g24_23, p24_23, g25_23, p25_23);
GREY grey25(g25_23, p25_23, g22_0, c25);
BLACK black24_23(g24_24, p24_24, g23_23, p23_23, g24_23, p24_23);
GREY grey24(g24_23, p24_23, g22_0, c24);
GREY grey23(g23_23, p23_23, g22_0, c23);
GREY grey22(g22_22, p22_22, g21_0, c22);
GREY grey21(g21_21, p21_21, g20_0, c21);
GREY grey20(g20_20, p20_20, g19_0, c20);
GREY grey19(g19_19, p19_19, g18_0, c19);
GREY grey18(g18_18, p18_18, g17_0, c18);
GREY grey17(g17_17, p17_17, g16_0, c17);
GREY grey16(g16_16, p16_16, g15_0, c16);
BLACK black15_8(g15_15, p15_15, g14_8, p14_8, g15_8, p15_8);
GREY grey15(g15_8, p15_8, g7_0, c15);
BLACK black14_8(g14_14, p14_14, g13_8, p13_8, g14_8, p14_8);
GREY grey14(g14_8, p14_8, g7_0, c14);
BLACK black13_8(g13_13, p13_13, g12_8, p12_8, g13_8, p13_8);
GREY grey13(g13_8, p13_8, g7_0, c13);
BLACK black12_8(g12_12, p12_12, g11_8, p11_8, g12_8, p12_8);
GREY grey12(g12_8, p12_8, g7_0, c12);
BLACK black11_8(g11_11, p11_11, g10_8, p10_8, g11_8, p11_8);
GREY grey11(g11_8, p11_8, g7_0, c11);
BLACK black10_8(g10_10, p10_10, g9_8, p9_8, g10_8, p10_8);
GREY grey10(g10_8, p10_8, g7_0, c10);
BLACK black9_8(g9_9, p9_9, g8_8, p8_8, g9_8, p9_8);
BLACK black9_7(g9_8, p9_8, g7_7, p7_7, g9_7, p9_7);
GREY grey9(g9_7, p9_7, g6_0, c9);
GREY grey8(g8_8, p8_8, g7_0, c8);
GREY grey7(g7_7, p7_7, g6_0, c7);
GREY grey6(g6_6, p6_6, g5_0, c6);
GREY grey5(g5_5, p5_5, g4_0, c5);
GREY grey4(g4_4, p4_4, g3_0, c4);
GREY grey3(g3_3, p3_3, g2_0, c3);
GREY grey2(g2_2, p2_2, g1_0, c2);
GREY grey1(g1_1, p1_1, g0_0, c1);
assign s[0] = a[0] ^ b[0];
assign c0 = g0_0;
assign cout = c63;
assign s[1] = p1_1 ^ c0;
assign s[2] = p2_2 ^ c1;
assign s[3] = p3_3 ^ c2;
assign s[4] = p4_4 ^ c3;
assign s[5] = p5_5 ^ c4;
assign s[6] = p6_6 ^ c5;
assign s[7] = p7_7 ^ c6;
assign s[8] = p8_8 ^ c7;
assign s[9] = p9_9 ^ c8;
assign s[10] = p10_10 ^ c9;
assign s[11] = p11_11 ^ c10;
assign s[12] = p12_12 ^ c11;
assign s[13] = p13_13 ^ c12;
assign s[14] = p14_14 ^ c13;
assign s[15] = p15_15 ^ c14;
assign s[16] = p16_16 ^ c15;
assign s[17] = p17_17 ^ c16;
assign s[18] = p18_18 ^ c17;
assign s[19] = p19_19 ^ c18;
assign s[20] = p20_20 ^ c19;
assign s[21] = p21_21 ^ c20;
assign s[22] = p22_22 ^ c21;
assign s[23] = p23_23 ^ c22;
assign s[24] = p24_24 ^ c23;
assign s[25] = p25_25 ^ c24;
assign s[26] = p26_26 ^ c25;
assign s[27] = p27_27 ^ c26;
assign s[28] = p28_28 ^ c27;
assign s[29] = p29_29 ^ c28;
assign s[30] = p30_30 ^ c29;
assign s[31] = p31_31 ^ c30;
assign s[32] = p32_32 ^ c31;
assign s[33] = p33_33 ^ c32;
assign s[34] = p34_34 ^ c33;
assign s[35] = p35_35 ^ c34;
assign s[36] = p36_36 ^ c35;
assign s[37] = p37_37 ^ c36;
assign s[38] = p38_38 ^ c37;
assign s[39] = p39_39 ^ c38;
assign s[40] = p40_40 ^ c39;
assign s[41] = p41_41 ^ c40;
assign s[42] = p42_42 ^ c41;
assign s[43] = p43_43 ^ c42;
assign s[44] = p44_44 ^ c43;
assign s[45] = p45_45 ^ c44;
assign s[46] = p46_46 ^ c45;
assign s[47] = p47_47 ^ c46;
assign s[48] = p48_48 ^ c47;
assign s[49] = p49_49 ^ c48;
assign s[50] = p50_50 ^ c49;
assign s[51] = p51_51 ^ c50;
assign s[52] = p52_52 ^ c51;
assign s[53] = p53_53 ^ c52;
assign s[54] = p54_54 ^ c53;
assign s[55] = p55_55 ^ c54;
assign s[56] = p56_56 ^ c55;
assign s[57] = p57_57 ^ c56;
assign s[58] = p58_58 ^ c57;
assign s[59] = p59_59 ^ c58;
assign s[60] = p60_60 ^ c59;
assign s[61] = p61_61 ^ c60;
assign s[62] = p62_62 ^ c61;
assign s[63] = p63_63 ^ c62;
endmodule

module GREY(gik, pik, gkj, gij);
input gik, pik, gkj;
output gij;
assign gij = gik | (pik & gkj);
endmodule

module BLACK(gik, pik, gkj, pkj, gij, pij);
input gik, pik, gkj, pkj;
output gij, pij;
assign pij = pik & pkj;
assign gij = gik | (pik & gkj);
endmodule

